.SUBCKT ASYNC_DFFHx1_ASAP7_75t_R CLK D QN RESET SET VDD VSS
MM43 pd3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM34 SH clkn pd3 VSS nmos_rvt w=81.0n l=20n nfin=3
MM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MM33 pd3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
MM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM37 pd2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MM35 SH clkb pd2 VDD pmos_rvt w=162.0n l=20n nfin=6
MM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M43 pd3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M34 SH clkn pd3 VSS nmos_rvt w=81.0n l=20n nfin=3
M48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
M33 pd3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
M8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
M47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
M25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
M22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M37 pd2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
M35 SH clkb pd2 VDD pmos_rvt w=162.0n l=20n nfin=6
M49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
M11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
M10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
M7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
M42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
M1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
M3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM43 pd3 SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM24 QN SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM29 SS SH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM23 clkb clkn VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM20 clkn CLK VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM44 SS RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM34 SH clkn pd3 VSS nmos_rvt w=81.0n l=20n nfin=3
MMM48 net020 RESET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM12 MS clkb SH VSS nmos_rvt w=81.0n l=20n nfin=3
MMM33 pd3 SS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM9 MH clkb net020 VSS nmos_rvt w=81.0n l=20n nfin=3
MMM8 net020 MS VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM6 MS MH VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM5 pd1 D VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM4 MH clkn pd1 VSS nmos_rvt w=81.0n l=20n nfin=3
MMM47 MS SET VSS VSS nmos_rvt w=81.0n l=20n nfin=3
MMM25 QN SH VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM28 SS SH net076 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM22 clkb clkn VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM45 net076 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM46 net079 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM21 clkn CLK VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM37 pd2 SS net077 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM35 SH clkb pd2 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM49 net078 RESET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM13 MS clkn SH VDD pmos_rvt w=162.0n l=20n nfin=6
MMM11 net051 MS net078 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM10 MH clkn net051 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM7 MS MH net079 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM42 net077 SET VDD VDD pmos_rvt w=162.0n l=20n nfin=6
MMM1 MH clkb pu1 VDD pmos_rvt w=162.0n l=20n nfin=6
MMM3 pu1 D VDD VDD pmos_rvt w=162.0n l=20n nfin=6
.ENDS